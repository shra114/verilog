/////////////////////////////////////////
//Description
// 
/////////////////////////////////////////
//import top_pkg::*;

module top (
  input  logic        clk,
  input  logic        rst_n 

);

//Internal signals

/////////////////////////
//Combinational logic
/////////////////////////

/////////////////////////
//Sequential logic
/////////////////////////
 
/////////////////////////
//Sub block instantiations
/////////////////////////

/////////////////////////
//Assertions
/////////////////////////
endmodule 
